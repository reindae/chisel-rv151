module control(
  input         clock,
  input         reset,
  input  [31:0] io_curr_inst,
  input  [31:0] io_prev_inst,
  input         io_BrEq,
  input         io_BrLt,
  input  [1:0]  io_curr_ALU_low2,
  input  [1:0]  io_prev_ALU_low2,
  output        io_PCSel,
  output [3:0]  io_ALUSel,
  output        io_BrUn,
  output        io_ASel,
  output        io_BSel,
  output        io_CSRSel,
  output        io_CSRWEn,
  output [31:0] io_DMEM_in,
  output [3:0]  io_DMEM_WEn,
  output [3:0]  io_DMEM_out,
  output        io_sign_ext,
  output [1:0]  io_WBSel,
  output        io_RegWEn,
  output        io_has_rd
);
  wire [6:0] curr_opc = io_curr_inst[6:0]; // @[control.scala 40:30]
  wire [2:0] curr_fn3 = io_curr_inst[14:12]; // @[control.scala 41:30]
  wire [6:0] prev_opc = io_prev_inst[6:0]; // @[control.scala 44:30]
  wire [2:0] prev_fn3 = io_prev_inst[14:12]; // @[control.scala 45:30]
  wire  _io_ALUSel_T_1 = ~io_curr_inst[30]; // @[control.scala 73:53]
  wire [3:0] _io_ALUSel_T_2 = ~io_curr_inst[30] ? 4'ha : 4'h6; // @[control.scala 73:34]
  wire [3:0] _io_ALUSel_T_4 = 3'h6 == curr_fn3 ? 4'h3 : 4'h1; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_6 = 3'h7 == curr_fn3 ? 4'h2 : _io_ALUSel_T_4; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_8 = 3'h4 == curr_fn3 ? 4'h4 : _io_ALUSel_T_6; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_10 = 3'h1 == curr_fn3 ? 4'h7 : _io_ALUSel_T_8; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_12 = 3'h2 == curr_fn3 ? 4'h8 : _io_ALUSel_T_10; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_14 = 3'h3 == curr_fn3 ? 4'h9 : _io_ALUSel_T_12; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_16 = 3'h5 == curr_fn3 ? _io_ALUSel_T_2 : _io_ALUSel_T_14; // @[Mux.scala 81:58]
  wire [6:0] _io_DMEM_WEn_T = 7'h1 << io_curr_ALU_low2; // @[control.scala 86:42]
  wire [1:0] _io_DMEM_WEn_T_2 = {1'h0,io_curr_ALU_low2[1]}; // @[Cat.scala 33:92]
  wire [2:0] _io_DMEM_WEn_T_3 = {_io_DMEM_WEn_T_2, 1'h0}; // @[control.scala 87:81]
  wire [10:0] _io_DMEM_WEn_T_4 = 11'h3 << _io_DMEM_WEn_T_3; // @[control.scala 87:42]
  wire [6:0] _io_DMEM_WEn_T_6 = 3'h0 == curr_fn3 ? _io_DMEM_WEn_T : 7'h0; // @[Mux.scala 81:58]
  wire [10:0] _io_DMEM_WEn_T_8 = 3'h1 == curr_fn3 ? _io_DMEM_WEn_T_4 : {{4'd0}, _io_DMEM_WEn_T_6}; // @[Mux.scala 81:58]
  wire [10:0] _io_DMEM_WEn_T_10 = 3'h2 == curr_fn3 ? 11'hf : _io_DMEM_WEn_T_8; // @[Mux.scala 81:58]
  wire [31:0] _io_DMEM_in_T_3 = 3'h0 == curr_fn3 ? 32'h1 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_DMEM_in_T_5 = 3'h1 == curr_fn3 ? 32'h1 : _io_DMEM_in_T_3; // @[Mux.scala 81:58]
  wire [31:0] _io_DMEM_in_T_7 = 3'h2 == curr_fn3 ? 32'h1 : _io_DMEM_in_T_5; // @[Mux.scala 81:58]
  wire  _io_PCSel_T = ~io_BrEq; // @[control.scala 103:27]
  wire  _io_PCSel_T_1 = ~io_BrLt; // @[control.scala 105:27]
  wire  _io_PCSel_T_6 = 3'h1 == curr_fn3 ? _io_PCSel_T : 3'h0 == curr_fn3 & io_BrEq; // @[Mux.scala 81:58]
  wire  _io_PCSel_T_8 = 3'h4 == curr_fn3 ? io_BrLt : _io_PCSel_T_6; // @[Mux.scala 81:58]
  wire  _io_PCSel_T_10 = 3'h5 == curr_fn3 ? _io_PCSel_T_1 : _io_PCSel_T_8; // @[Mux.scala 81:58]
  wire  _io_PCSel_T_12 = 3'h6 == curr_fn3 ? io_BrLt : _io_PCSel_T_10; // @[Mux.scala 81:58]
  wire  _io_PCSel_T_14 = 3'h7 == curr_fn3 ? _io_PCSel_T_1 : _io_PCSel_T_12; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_19 = _io_ALUSel_T_1 ? 4'h1 : 4'h5; // @[control.scala 145:35]
  wire [3:0] _io_ALUSel_T_24 = 3'h6 == curr_fn3 ? 4'h3 : _io_ALUSel_T_19; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_26 = 3'h7 == curr_fn3 ? 4'h2 : _io_ALUSel_T_24; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_28 = 3'h4 == curr_fn3 ? 4'h4 : _io_ALUSel_T_26; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_30 = 3'h1 == curr_fn3 ? 4'h7 : _io_ALUSel_T_28; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_32 = 3'h2 == curr_fn3 ? 4'h8 : _io_ALUSel_T_30; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_34 = 3'h3 == curr_fn3 ? 4'h9 : _io_ALUSel_T_32; // @[Mux.scala 81:58]
  wire [3:0] _io_ALUSel_T_36 = 3'h5 == curr_fn3 ? _io_ALUSel_T_2 : _io_ALUSel_T_34; // @[Mux.scala 81:58]
  wire [3:0] _GEN_0 = 7'h33 == curr_opc ? _io_ALUSel_T_36 : 4'h0; // @[control.scala 144:17 48:13 62:21]
  wire  _GEN_1 = 7'h73 == curr_opc & curr_fn3 == 3'h5; // @[control.scala 139:17 53:13 62:21]
  wire [3:0] _GEN_3 = 7'h73 == curr_opc ? 4'h0 : _GEN_0; // @[control.scala 48:13 62:21]
  wire [3:0] _GEN_5 = 7'h37 == curr_opc ? 4'hb : _GEN_3; // @[control.scala 135:17 62:21]
  wire  _GEN_6 = 7'h37 == curr_opc ? 1'h0 : _GEN_1; // @[control.scala 53:13 62:21]
  wire  _GEN_7 = 7'h37 == curr_opc ? 1'h0 : 7'h73 == curr_opc; // @[control.scala 52:13 62:21]
  wire  _GEN_8 = 7'h17 == curr_opc | 7'h37 == curr_opc; // @[control.scala 127:15 62:21]
  wire [3:0] _GEN_9 = 7'h17 == curr_opc ? 4'h1 : _GEN_5; // @[control.scala 129:17 62:21]
  wire  _GEN_10 = 7'h17 == curr_opc ? 1'h0 : _GEN_6; // @[control.scala 53:13 62:21]
  wire  _GEN_11 = 7'h17 == curr_opc ? 1'h0 : _GEN_7; // @[control.scala 52:13 62:21]
  wire  _GEN_13 = 7'h67 == curr_opc ? 1'h0 : _GEN_8; // @[control.scala 121:15 62:21]
  wire  _GEN_14 = 7'h67 == curr_opc | _GEN_8; // @[control.scala 122:15 62:21]
  wire [3:0] _GEN_15 = 7'h67 == curr_opc ? 4'h1 : _GEN_9; // @[control.scala 123:17 62:21]
  wire  _GEN_16 = 7'h67 == curr_opc ? 1'h0 : _GEN_10; // @[control.scala 53:13 62:21]
  wire  _GEN_17 = 7'h67 == curr_opc ? 1'h0 : _GEN_11; // @[control.scala 52:13 62:21]
  wire  _GEN_18 = 7'h6f == curr_opc | 7'h67 == curr_opc; // @[control.scala 113:16 62:21]
  wire  _GEN_19 = 7'h6f == curr_opc | _GEN_13; // @[control.scala 114:15 62:21]
  wire  _GEN_20 = 7'h6f == curr_opc | _GEN_14; // @[control.scala 115:15 62:21]
  wire [3:0] _GEN_21 = 7'h6f == curr_opc ? 4'h1 : _GEN_15; // @[control.scala 116:17 62:21]
  wire  _GEN_22 = 7'h6f == curr_opc ? 1'h0 : _GEN_16; // @[control.scala 53:13 62:21]
  wire  _GEN_23 = 7'h6f == curr_opc ? 1'h0 : _GEN_17; // @[control.scala 52:13 62:21]
  wire  _GEN_24 = 7'h63 == curr_opc | _GEN_19; // @[control.scala 62:21 98:15]
  wire  _GEN_25 = 7'h63 == curr_opc | _GEN_20; // @[control.scala 62:21 99:15]
  wire [3:0] _GEN_26 = 7'h63 == curr_opc ? 4'h1 : _GEN_21; // @[control.scala 100:17 62:21]
  wire  _GEN_27 = 7'h63 == curr_opc ? _io_PCSel_T_14 : _GEN_18; // @[control.scala 101:16 62:21]
  wire  _GEN_28 = 7'h63 == curr_opc & (curr_fn3 == 3'h6 | curr_fn3 == 3'h7); // @[control.scala 109:15 49:11 62:21]
  wire  _GEN_29 = 7'h63 == curr_opc ? 1'h0 : _GEN_22; // @[control.scala 53:13 62:21]
  wire  _GEN_30 = 7'h63 == curr_opc ? 1'h0 : _GEN_23; // @[control.scala 52:13 62:21]
  wire  _GEN_31 = 7'h23 == curr_opc | _GEN_25; // @[control.scala 62:21 83:15]
  wire [3:0] _GEN_32 = 7'h23 == curr_opc ? 4'h1 : _GEN_26; // @[control.scala 62:21 84:17]
  wire [10:0] _GEN_33 = 7'h23 == curr_opc ? _io_DMEM_WEn_T_10 : 11'h0; // @[control.scala 54:15 62:21 85:19]
  wire [31:0] _GEN_34 = 7'h23 == curr_opc ? _io_DMEM_in_T_7 : 32'h0; // @[control.scala 55:14 62:21 90:18]
  wire  _GEN_35 = 7'h23 == curr_opc ? 1'h0 : _GEN_24; // @[control.scala 50:11 62:21]
  wire  _GEN_36 = 7'h23 == curr_opc ? 1'h0 : _GEN_27; // @[control.scala 47:12 62:21]
  wire  _GEN_37 = 7'h23 == curr_opc ? 1'h0 : _GEN_28; // @[control.scala 49:11 62:21]
  wire  _GEN_38 = 7'h23 == curr_opc ? 1'h0 : _GEN_29; // @[control.scala 53:13 62:21]
  wire  _GEN_39 = 7'h23 == curr_opc ? 1'h0 : _GEN_30; // @[control.scala 52:13 62:21]
  wire  _GEN_40 = 7'h3 == curr_opc | _GEN_31; // @[control.scala 62:21 78:15]
  wire [3:0] _GEN_41 = 7'h3 == curr_opc ? 4'h1 : _GEN_32; // @[control.scala 62:21 79:17]
  wire [10:0] _GEN_42 = 7'h3 == curr_opc ? 11'h0 : _GEN_33; // @[control.scala 54:15 62:21]
  wire [31:0] _GEN_43 = 7'h3 == curr_opc ? 32'h0 : _GEN_34; // @[control.scala 55:14 62:21]
  wire  _GEN_44 = 7'h3 == curr_opc ? 1'h0 : _GEN_35; // @[control.scala 50:11 62:21]
  wire  _GEN_45 = 7'h3 == curr_opc ? 1'h0 : _GEN_36; // @[control.scala 47:12 62:21]
  wire  _GEN_46 = 7'h3 == curr_opc ? 1'h0 : _GEN_37; // @[control.scala 49:11 62:21]
  wire  _GEN_47 = 7'h3 == curr_opc ? 1'h0 : _GEN_38; // @[control.scala 53:13 62:21]
  wire  _GEN_48 = 7'h3 == curr_opc ? 1'h0 : _GEN_39; // @[control.scala 52:13 62:21]
  wire [10:0] _GEN_51 = 7'h13 == curr_opc ? 11'h0 : _GEN_42; // @[control.scala 54:15 62:21]
  wire  _io_RegWEn_T_1 = io_prev_inst[11:7] != 5'h0; // @[control.scala 159:39]
  wire  _io_sign_ext_T_3 = prev_fn3 == 3'h4 | prev_fn3 == 3'h5 ? 1'h0 : 1'h1; // @[control.scala 172:25]
  wire [1:0] _io_DMEM_out_T_1 = {1'h0,io_prev_ALU_low2[1]}; // @[Cat.scala 33:92]
  wire [2:0] _io_DMEM_out_T_2 = {_io_DMEM_out_T_1, 1'h0}; // @[control.scala 175:81]
  wire [10:0] _io_DMEM_out_T_3 = 11'h3 << _io_DMEM_out_T_2; // @[control.scala 175:42]
  wire [6:0] _io_DMEM_out_T_8 = 7'h1 << io_prev_ALU_low2; // @[control.scala 177:42]
  wire [3:0] _io_DMEM_out_T_11 = 3'h2 == prev_fn3 ? 4'hf : 4'h0; // @[Mux.scala 81:58]
  wire [10:0] _io_DMEM_out_T_13 = 3'h2 == prev_fn3 ? _io_DMEM_out_T_3 : {{7'd0}, _io_DMEM_out_T_11}; // @[Mux.scala 81:58]
  wire [10:0] _io_DMEM_out_T_15 = 3'h2 == prev_fn3 ? _io_DMEM_out_T_3 : _io_DMEM_out_T_13; // @[Mux.scala 81:58]
  wire [10:0] _io_DMEM_out_T_17 = 3'h2 == prev_fn3 ? {{4'd0}, _io_DMEM_out_T_8} : _io_DMEM_out_T_15; // @[Mux.scala 81:58]
  wire [10:0] _io_DMEM_out_T_19 = 3'h2 == prev_fn3 ? {{4'd0}, _io_DMEM_out_T_8} : _io_DMEM_out_T_17; // @[Mux.scala 81:58]
  wire  _GEN_58 = 7'h73 == prev_opc & _io_RegWEn_T_1; // @[control.scala 157:21 183:17 60:13]
  wire  _GEN_59 = 7'h3 == prev_opc & _io_RegWEn_T_1; // @[control.scala 157:21 171:17 59:13]
  wire  _GEN_60 = 7'h3 == prev_opc & _io_sign_ext_T_3; // @[control.scala 157:21 172:19 57:15]
  wire [10:0] _GEN_61 = 7'h3 == prev_opc ? _io_DMEM_out_T_19 : 11'h0; // @[control.scala 157:21 173:19 56:15]
  wire  _GEN_62 = 7'h3 == prev_opc ? 1'h0 : _GEN_58; // @[control.scala 157:21 60:13]
  wire  _GEN_63 = 7'h6f == prev_opc | 7'h67 == prev_opc ? _io_RegWEn_T_1 : _GEN_59; // @[control.scala 157:21 165:17]
  wire [1:0] _GEN_64 = 7'h6f == prev_opc | 7'h67 == prev_opc ? 2'h2 : 2'h0; // @[control.scala 157:21 166:16 58:12]
  wire  _GEN_65 = 7'h6f == prev_opc | 7'h67 == prev_opc ? _io_RegWEn_T_1 : _GEN_62; // @[control.scala 157:21 167:17]
  wire  _GEN_66 = 7'h6f == prev_opc | 7'h67 == prev_opc ? 1'h0 : _GEN_60; // @[control.scala 157:21 57:15]
  wire [10:0] _GEN_67 = 7'h6f == prev_opc | 7'h67 == prev_opc ? 11'h0 : _GEN_61; // @[control.scala 157:21 56:15]
  wire [10:0] _GEN_72 = 7'h33 == prev_opc | 7'h13 == prev_opc | 7'h17 == prev_opc | 7'h37 == prev_opc ? 11'h0 : _GEN_67; // @[control.scala 157:21 56:15]
  assign io_PCSel = 7'h13 == curr_opc ? 1'h0 : _GEN_45; // @[control.scala 47:12 62:21]
  assign io_ALUSel = 7'h13 == curr_opc ? _io_ALUSel_T_16 : _GEN_41; // @[control.scala 62:21 65:17]
  assign io_BrUn = 7'h13 == curr_opc ? 1'h0 : _GEN_46; // @[control.scala 49:11 62:21]
  assign io_ASel = 7'h13 == curr_opc ? 1'h0 : _GEN_44; // @[control.scala 50:11 62:21]
  assign io_BSel = 7'h13 == curr_opc | _GEN_40; // @[control.scala 62:21 64:15]
  assign io_CSRSel = 7'h13 == curr_opc ? 1'h0 : _GEN_47; // @[control.scala 53:13 62:21]
  assign io_CSRWEn = 7'h13 == curr_opc ? 1'h0 : _GEN_48; // @[control.scala 52:13 62:21]
  assign io_DMEM_in = 7'h13 == curr_opc ? 32'h0 : _GEN_43; // @[control.scala 55:14 62:21]
  assign io_DMEM_WEn = _GEN_51[3:0];
  assign io_DMEM_out = _GEN_72[3:0];
  assign io_sign_ext = 7'h33 == prev_opc | 7'h13 == prev_opc | 7'h17 == prev_opc | 7'h37 == prev_opc ? 1'h0 : _GEN_66; // @[control.scala 157:21 57:15]
  assign io_WBSel = 7'h33 == prev_opc | 7'h13 == prev_opc | 7'h17 == prev_opc | 7'h37 == prev_opc ? 2'h1 : _GEN_64; // @[control.scala 157:21 160:16]
  assign io_RegWEn = 7'h33 == prev_opc | 7'h13 == prev_opc | 7'h17 == prev_opc | 7'h37 == prev_opc ? io_prev_inst[11:7]
     != 5'h0 : _GEN_63; // @[control.scala 157:21 159:17]
  assign io_has_rd = 7'h33 == prev_opc | 7'h13 == prev_opc | 7'h17 == prev_opc | 7'h37 == prev_opc ? _io_RegWEn_T_1 :
    _GEN_65; // @[control.scala 157:21 161:17]
endmodule
